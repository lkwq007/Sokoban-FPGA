library verilog;
use verilog.vl_types.all;
entity game_core_tb is
    generic(
        DELAY           : integer := 100
    );
end game_core_tb;
