library verilog;
use verilog.vl_types.all;
entity ms_gen_lfsr_tb is
end ms_gen_lfsr_tb;
