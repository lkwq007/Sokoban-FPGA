library verilog;
use verilog.vl_types.all;
entity ps2_dataprogramme_tb is
end ps2_dataprogramme_tb;
