library verilog;
use verilog.vl_types.all;
entity game_controller_tb is
    generic(
        DELAY           : integer := 10
    );
end game_controller_tb;
