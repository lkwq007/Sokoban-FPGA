library verilog;
use verilog.vl_types.all;
entity ms_gen_tb is
end ms_gen_tb;
