library verilog;
use verilog.vl_types.all;
entity ms_controller_tb is
end ms_controller_tb;
