library verilog;
use verilog.vl_types.all;
entity svga_top_tb is
end svga_top_tb;
