library verilog;
use verilog.vl_types.all;
entity game_man_move_tb is
    generic(
        DELAY           : integer := 10
    );
end game_man_move_tb;
