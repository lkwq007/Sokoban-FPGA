library verilog;
use verilog.vl_types.all;
entity mouse_interterface_tb_v is
end mouse_interterface_tb_v;
