library verilog;
use verilog.vl_types.all;
entity ms_round_tb is
end ms_round_tb;
